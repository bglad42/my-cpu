`timescale 1ns/1ps
module pipelined (clk, reset);
	input logic clk, reset;
	wire notClk
	// generate instruction!
	
	wire [31:0] instr_toreg, instr;
	wire [63:0] pc, newpc;
	logic UncondBr, BrTaken, Reg2Loc, RegWrite, MemWrite, MemToReg; // controls
	logic [2:0] ALUOp; // more control
	logic [1:0] ALUSrc; // more
	
	// flags
	
	logic zero, overflow, carryout, negative, flagWrite;
	wire ALUz, ALUo, ALUc, ALUn;
	
	D_FF_en zeroFlag 		(.q(zero), 		.d(ALUz), .clk(clk), .reset(reset), .en(flagWrite));
	D_FF_en overflowFlag (.q(overflow), .d(ALUo), .clk(clk), .reset(reset), .en(flagWrite));
	D_FF_en carryoutFlag (.q(carryout), .d(ALUc), .clk(clk), .reset(reset), .en(flagWrite));
	D_FF_en negativeFlag (.q(negative), .d(ALUn), .clk(clk), .reset(reset), .en(flagWrite));
	
	
	//  Instruction fetch (IF)
	// ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
	
	programCounter current (.q(pc), .d(newpc), .clk(clk), .reset(reset)); // out to pc, in from newpc
	
	instructmem instruction (.instruction(instr), .address(pc), .clk(clk));
	
	// ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
	
	
	IF_ID IF_ID_register (.PCin(), .PCout(), .instr(instr_toreg), instr_out(instr), .clk, .reset); // finish via last pipeline register
	
	
	// Register Fetch (ID)
	// ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
	
	logic [4:0] Rd, Rm, Rn;
	assign Rd = instr[4:0];
	assign Rn = instr[9:5];
	assign Rm = instr[20:16];
	
	wire [63:0] Dw, Da, Db;
	wire [4:0] Bin;
						
	wire [63:0] ALUResult, DAddr, ALUBin, Imm, LSR;
	
	sign_extend #(.WIDTH(9)) Addr (.out(DAddr), .in(instr[20:12]));
	zero_extend #(.WIDTH(12)) Imm12 (.out(Imm), .in(instr[21:10]));
	
	shifter LogicalShiftRight (.value(Da), .direction(1'b1), .distance(instr[15:10]), .result(LSR));
	
	generate
		for (i = 0; i < 64; i++) begin : each4Mux
			wire [3:0] temp;
			assign temp[0] = Db[i];
			assign temp[1] = DAddr[i];
			assign temp[2] = Imm[i];
			assign temp[3] = LSR[i];
			mux4_1 alusourcer (.out(ALUBin[i]), .in(temp), .sel(ALUSrc));
		end
	endgenerate
	
	not #50 clkHack (notClk, clk);
	
	regfile reggie (.ReadData1(Da), .ReadData2(Db), .WriteData(Dw), .ReadRegister1(Rn),
						.ReadRegister2(Bin), .WriteRegister(Rd), .RegWrite(RegWrite), .clk(notClk), .reset);
	
	controls broisthethinker (.Reg2Loc(Reg2Loc), .UncondBr(UncondBr), .BrTaken(BrTaken), .RegWrite(RegWrite), 
									  .MemWrite(MemWrite), .ALUOp(ALUOp), .ALUSrc(ALUSrc), .MemToReg(MemToReg), 
									  .instr(instr), .zero(zero), .negative(negative), .overflow(overflow), 
									  .flagWrite(flagWrite), .ALUz(ALUz));
	// end register fetch
	// ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~					
						
						
	ID_EX ID_EX_register (.RegWrite(), .MemWrite(), .ALUOp(), .ALUSrc(), .MemToReg(), .flagWrite(), 
								.RegWrite_out(), .MemWrite_out(), .ALUOp_out(), .ALUSrc_out(), .MemToReg_out(), .instr_out(), .flagWrite_out(),
								.Imm12Ext(), .Daddr9Ext(), .LS(), .Rd(), .Da(), .Db(), .Imm12Ext_out(), .Daddr9Ext_out(), .LS_out(), .Rd_out(),
								.Da_out(), .Db_out(), .clk, .reset);
								
	// Execute (EX)
	// ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
	
		alu ALU (.result(ALUResult), .A(Da), .B(ALUBin), .cntrl(ALUOp), .negative(ALUn), .zero(ALUz), .overflow(ALUo), .carry_out(ALUc)); //might need flag registers?

	// ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
	
	
	EX_MEM EX_MEM_register (.Db(), .Daddr9Ext(), .MemWrite(), .MemToReg(), .FlagWrite(), .RegWrite(), .Rd(), .clk, .reset, 
									.Db_out(), .Daddr9Ext_out(), .MemWrite_out(), .MemToReg_out(), .FlagWrite_out(), .RegWrite_out(), .Rd_out());
	

	// Data Memory (MEM)
	// ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
	
	wire [63:0] memDataOut;
	datamem dataMemory (.address(ALUResult), .write_enable(MemWrite), .read_enable(1'b1), // read up on xfer size, read enable reqs
								.write_data(Db), .clk(clk), .xfer_size(4'b1000), .read_data(memDataOut));
	
	// ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
	
	
	MEM_WR MEM_WR_register (.RegWrite(), .RegWrite_out(), .Rd(), .Rd_out(), .Data(), .DataOut(), .clk, .reset);
	
	
	// Writeback (WR)
	// ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
	
	mux_64_2_1 toReg (.out(Dw), .A(ALUResult), .B(memDataOut), .sel(MemToReg));
	
	// ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~

	
	wire [63:0] updateloc, uncond, cond, branch, nobranch, branchPC;
	
	sign_extend #(.WIDTH(26)) unc (.out(uncond), .in(instr[25:0])); // se BrAddr26
	sign_extend #(.WIDTH(19)) con (.out(cond), .in(instr[23:5])); // se CondAddr19
	
	mux_64_2_1 CondUncond (.out(updateloc), .A(cond), .B(uncond), .sel(UncondBr)); // selecting UncondBranch or not
	
	shifter shifty (.value(updateloc), .direction(1'b0), .distance(6'd2), .result(branch)); //shift result 2 for branch addition
	
	adder_64 BranchPCUpdate (.out(branchPC), .A(pc), .B(branch)); // add branch to pc, send to branchPC for update
	adder_64 PCUpdate (.out(nobranch), .A(pc), .B(64'd4)); // update pc on no branch
	mux_64_2_1 branchOrNot (.out(newpc), .A(nobranch), .B(branchPC), .sel(BrTaken)); // select new pc address 
	
	
endmodule

module pipelined_testbench();
	
	logic clk, reset;
	
	parameter ClockDelay = 20000;
	pipelined dut (.clk(clk), .reset(reset));
	
	initial begin // Set up the clock
		clk <= 0;
		forever #(ClockDelay/2) clk <= ~clk;
	end
	
	int i;
	initial begin
		reset = 1;	@(posedge clk);
		reset = 0;	@(posedge clk);
		for (i = 0; i < 100; i++) begin
			@(posedge clk);
		end
		$stop;
	end
endmodule