module ID_EX (//controls
					RegWrite, MemWrite, ALUOp, ALUSrc, MemToReg, flagWrite, 
					RegWrite_out, MemWrite_out, ALUOp_out, ALUSrc_out, MemToReg_out, instr_out, flagWrite_out
					// operations/operators
					Imm12Ext, Daddr9Ext, LS, Rd, Da, Db,
					Imm12Ext_out, Daddr9Ext_out, LS_out, Rd_out, Da_out, Db_out,
					// inputs
					clk, reset);
	
	input logic RegWrite, MemWrite, MemToReg, flagWrite, clk, reset;
	input logic [1:0] ALUSrc;
	input logic [2:0] ALUOp;
	input logic [4:0] Rd;
	input logic [63:0] Da, Db, LS; 
	output logic RegWrite_out, MemWrite_out, ALUOp_out, ALUSrc_out, MemToReg_out, instr_out, flagWrite_out;
	output logic [1:0] ALUSrc_out;
	output logic [2:0] ALUOp_out;
	output logic [4:0] Rd_out;
	output logic [63:0] Da_out, Db_out, LS_out;
					
	
	D_FF RegWriteID (.q(RegWrite_out), .d(RegWrite), .clk, .reset);
	D_FF MemWriteID (.q(MemWrite_out), .d(MemWrite), .clk, .reset);
	D_FF FlagWriteID (.q(flagWrite_out), .d(flagWrite), .clk, .reset);
	
	regmodular #(.WIDTH(2)) ALUSrcReg (.out(ALUSrc_out), .in(ALUSrc), .clk, .reset);
	regmodular #(.WIDTH(3)) ALUOpReg (.out(ALUOp_out), .in(ALUOp), .clk, .reset);
	regmodular #(.WIDTH(64)) DaReg (.out(Da_out), .in(Da), .clk, .reset);
	regmodular #(.WIDTH(64)) DbReg (.out(Db_out), .in(Db), .clk, .reset);
endmodule 